library verilog;
use verilog.vl_types.all;
entity beep_tb is
end beep_tb;
